module simple_logic (input a, b, output y); assign y = a & b; endmodule
