module complex_logic (input x, y, z, output w); assign w = (x & y) | z; endmodule
